module fifo(
    input rst,
    input wr_clk,
    input wr_en,
    input [7:0] din,

    input rd_clk,
    input rd_en,
    output [7:0] dout
);



endmodule