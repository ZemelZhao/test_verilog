module cs_cmd(
    input clk,
    input rst,
);

    

endmodule