module cs_clk(
    input clk,
    output spi_clk,
    output fs_adc
);
    
    

endmodule