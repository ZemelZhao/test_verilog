module cs_cmd(
    input sys_clk,
    input rst,

    input fs_adc,

    input fs_udp_rx,
    output fs_udp_tx,
    output fs_fifod2mac,
    output fs_mac2fifoc,
    output fs_fifoc2cs,
    output fs_adc_check,
    output fs_adc_conf,
    output fs_adc_read,
    output fs_adc_fifo,

    output fd_udp_rx,
    input fd_udp_tx,
    input fd_fifod2mac,
    input fd_mac2fifoc,
    input fd_fifoc2cs,
    input fd_adc_check,
    input fd_adc_conf,
    input fd_adc_read,
    input fd_adc_fifo
);

    




endmodule