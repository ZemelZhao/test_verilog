module cs_clk(

);
    

endmodule