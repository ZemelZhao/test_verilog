module cs(
    input clk,
    input rst,

    input fifoa_full,
    input fifoc_full,
    input fifod_full

    
);



endmodule